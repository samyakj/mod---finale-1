`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:32:07 06/21/2014 
// Design Name: 
// Module Name:    mew 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module mew(output reg[63:0] new
    );
new<=64'b10101010_10101010_10101010_10101010_10101010_10101010_10101010_10101010;

endmodule
